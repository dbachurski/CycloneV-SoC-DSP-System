/**
 * Copyright (C) 2023  AGH University of Science and Technology
 */

module and2 (
    output logic y,
    input logic  a,
    input logic  b
);


/**
 * Signals assignments
 */

assign y = a & b;

endmodule
